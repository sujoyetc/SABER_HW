`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:06:24 07/07/2019 
// Design Name: 
// Module Name:    parallel_Mults 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module parallel_Mults1(clk, acc, secret, a_coeff, result);
input clk;
input [3327:0] acc;
input [3327:0] secret;
input [12:0] a_coeff;
output [3327:0] result;

small_alu1 sa0(clk, acc[12:0], secret[12:0], a_coeff, result[12:0]);
small_alu1 sa1(clk, acc[25:13], secret[25:13], a_coeff, result[25:13]);
small_alu1 sa2(clk, acc[38:26], secret[38:26], a_coeff, result[38:26]);
small_alu1 sa3(clk, acc[51:39], secret[51:39], a_coeff, result[51:39]);
small_alu1 sa4(clk, acc[64:52], secret[64:52], a_coeff, result[64:52]);
small_alu1 sa5(clk, acc[77:65], secret[77:65], a_coeff, result[77:65]);
small_alu1 sa6(clk, acc[90:78], secret[90:78], a_coeff, result[90:78]);
small_alu1 sa7(clk, acc[103:91], secret[103:91], a_coeff, result[103:91]);
small_alu1 sa8(clk, acc[116:104], secret[116:104], a_coeff, result[116:104]);
small_alu1 sa9(clk, acc[129:117], secret[129:117], a_coeff, result[129:117]);
small_alu1 sa10(clk, acc[142:130], secret[142:130], a_coeff, result[142:130]);
small_alu1 sa11(clk, acc[155:143], secret[155:143], a_coeff, result[155:143]);
small_alu1 sa12(clk, acc[168:156], secret[168:156], a_coeff, result[168:156]);
small_alu1 sa13(clk, acc[181:169], secret[181:169], a_coeff, result[181:169]);
small_alu1 sa14(clk, acc[194:182], secret[194:182], a_coeff, result[194:182]);
small_alu1 sa15(clk, acc[207:195], secret[207:195], a_coeff, result[207:195]);
small_alu1 sa16(clk, acc[220:208], secret[220:208], a_coeff, result[220:208]);
small_alu1 sa17(clk, acc[233:221], secret[233:221], a_coeff, result[233:221]);
small_alu1 sa18(clk, acc[246:234], secret[246:234], a_coeff, result[246:234]);
small_alu1 sa19(clk, acc[259:247], secret[259:247], a_coeff, result[259:247]);
small_alu1 sa20(clk, acc[272:260], secret[272:260], a_coeff, result[272:260]);
small_alu1 sa21(clk, acc[285:273], secret[285:273], a_coeff, result[285:273]);
small_alu1 sa22(clk, acc[298:286], secret[298:286], a_coeff, result[298:286]);
small_alu1 sa23(clk, acc[311:299], secret[311:299], a_coeff, result[311:299]);
small_alu1 sa24(clk, acc[324:312], secret[324:312], a_coeff, result[324:312]);
small_alu1 sa25(clk, acc[337:325], secret[337:325], a_coeff, result[337:325]);
small_alu1 sa26(clk, acc[350:338], secret[350:338], a_coeff, result[350:338]);
small_alu1 sa27(clk, acc[363:351], secret[363:351], a_coeff, result[363:351]);
small_alu1 sa28(clk, acc[376:364], secret[376:364], a_coeff, result[376:364]);
small_alu1 sa29(clk, acc[389:377], secret[389:377], a_coeff, result[389:377]);
small_alu1 sa30(clk, acc[402:390], secret[402:390], a_coeff, result[402:390]);
small_alu1 sa31(clk, acc[415:403], secret[415:403], a_coeff, result[415:403]);
small_alu1 sa32(clk, acc[428:416], secret[428:416], a_coeff, result[428:416]);
small_alu1 sa33(clk, acc[441:429], secret[441:429], a_coeff, result[441:429]);
small_alu1 sa34(clk, acc[454:442], secret[454:442], a_coeff, result[454:442]);
small_alu1 sa35(clk, acc[467:455], secret[467:455], a_coeff, result[467:455]);
small_alu1 sa36(clk, acc[480:468], secret[480:468], a_coeff, result[480:468]);
small_alu1 sa37(clk, acc[493:481], secret[493:481], a_coeff, result[493:481]);
small_alu1 sa38(clk, acc[506:494], secret[506:494], a_coeff, result[506:494]);
small_alu1 sa39(clk, acc[519:507], secret[519:507], a_coeff, result[519:507]);
small_alu1 sa40(clk, acc[532:520], secret[532:520], a_coeff, result[532:520]);
small_alu1 sa41(clk, acc[545:533], secret[545:533], a_coeff, result[545:533]);
small_alu1 sa42(clk, acc[558:546], secret[558:546], a_coeff, result[558:546]);
small_alu1 sa43(clk, acc[571:559], secret[571:559], a_coeff, result[571:559]);
small_alu1 sa44(clk, acc[584:572], secret[584:572], a_coeff, result[584:572]);
small_alu1 sa45(clk, acc[597:585], secret[597:585], a_coeff, result[597:585]);
small_alu1 sa46(clk, acc[610:598], secret[610:598], a_coeff, result[610:598]);
small_alu1 sa47(clk, acc[623:611], secret[623:611], a_coeff, result[623:611]);
small_alu1 sa48(clk, acc[636:624], secret[636:624], a_coeff, result[636:624]);
small_alu1 sa49(clk, acc[649:637], secret[649:637], a_coeff, result[649:637]);
small_alu1 sa50(clk, acc[662:650], secret[662:650], a_coeff, result[662:650]);
small_alu1 sa51(clk, acc[675:663], secret[675:663], a_coeff, result[675:663]);
small_alu1 sa52(clk, acc[688:676], secret[688:676], a_coeff, result[688:676]);
small_alu1 sa53(clk, acc[701:689], secret[701:689], a_coeff, result[701:689]);
small_alu1 sa54(clk, acc[714:702], secret[714:702], a_coeff, result[714:702]);
small_alu1 sa55(clk, acc[727:715], secret[727:715], a_coeff, result[727:715]);
small_alu1 sa56(clk, acc[740:728], secret[740:728], a_coeff, result[740:728]);
small_alu1 sa57(clk, acc[753:741], secret[753:741], a_coeff, result[753:741]);
small_alu1 sa58(clk, acc[766:754], secret[766:754], a_coeff, result[766:754]);
small_alu1 sa59(clk, acc[779:767], secret[779:767], a_coeff, result[779:767]);
small_alu1 sa60(clk, acc[792:780], secret[792:780], a_coeff, result[792:780]);
small_alu1 sa61(clk, acc[805:793], secret[805:793], a_coeff, result[805:793]);
small_alu1 sa62(clk, acc[818:806], secret[818:806], a_coeff, result[818:806]);
small_alu1 sa63(clk, acc[831:819], secret[831:819], a_coeff, result[831:819]);
small_alu1 sa64(clk, acc[844:832], secret[844:832], a_coeff, result[844:832]);
small_alu1 sa65(clk, acc[857:845], secret[857:845], a_coeff, result[857:845]);
small_alu1 sa66(clk, acc[870:858], secret[870:858], a_coeff, result[870:858]);
small_alu1 sa67(clk, acc[883:871], secret[883:871], a_coeff, result[883:871]);
small_alu1 sa68(clk, acc[896:884], secret[896:884], a_coeff, result[896:884]);
small_alu1 sa69(clk, acc[909:897], secret[909:897], a_coeff, result[909:897]);
small_alu1 sa70(clk, acc[922:910], secret[922:910], a_coeff, result[922:910]);
small_alu1 sa71(clk, acc[935:923], secret[935:923], a_coeff, result[935:923]);
small_alu1 sa72(clk, acc[948:936], secret[948:936], a_coeff, result[948:936]);
small_alu1 sa73(clk, acc[961:949], secret[961:949], a_coeff, result[961:949]);
small_alu1 sa74(clk, acc[974:962], secret[974:962], a_coeff, result[974:962]);
small_alu1 sa75(clk, acc[987:975], secret[987:975], a_coeff, result[987:975]);
small_alu1 sa76(clk, acc[1000:988], secret[1000:988], a_coeff, result[1000:988]);
small_alu1 sa77(clk, acc[1013:1001], secret[1013:1001], a_coeff, result[1013:1001]);
small_alu1 sa78(clk, acc[1026:1014], secret[1026:1014], a_coeff, result[1026:1014]);
small_alu1 sa79(clk, acc[1039:1027], secret[1039:1027], a_coeff, result[1039:1027]);
small_alu1 sa80(clk, acc[1052:1040], secret[1052:1040], a_coeff, result[1052:1040]);
small_alu1 sa81(clk, acc[1065:1053], secret[1065:1053], a_coeff, result[1065:1053]);
small_alu1 sa82(clk, acc[1078:1066], secret[1078:1066], a_coeff, result[1078:1066]);
small_alu1 sa83(clk, acc[1091:1079], secret[1091:1079], a_coeff, result[1091:1079]);
small_alu1 sa84(clk, acc[1104:1092], secret[1104:1092], a_coeff, result[1104:1092]);
small_alu1 sa85(clk, acc[1117:1105], secret[1117:1105], a_coeff, result[1117:1105]);
small_alu1 sa86(clk, acc[1130:1118], secret[1130:1118], a_coeff, result[1130:1118]);
small_alu1 sa87(clk, acc[1143:1131], secret[1143:1131], a_coeff, result[1143:1131]);
small_alu1 sa88(clk, acc[1156:1144], secret[1156:1144], a_coeff, result[1156:1144]);
small_alu1 sa89(clk, acc[1169:1157], secret[1169:1157], a_coeff, result[1169:1157]);
small_alu1 sa90(clk, acc[1182:1170], secret[1182:1170], a_coeff, result[1182:1170]);
small_alu1 sa91(clk, acc[1195:1183], secret[1195:1183], a_coeff, result[1195:1183]);
small_alu1 sa92(clk, acc[1208:1196], secret[1208:1196], a_coeff, result[1208:1196]);
small_alu1 sa93(clk, acc[1221:1209], secret[1221:1209], a_coeff, result[1221:1209]);
small_alu1 sa94(clk, acc[1234:1222], secret[1234:1222], a_coeff, result[1234:1222]);
small_alu1 sa95(clk, acc[1247:1235], secret[1247:1235], a_coeff, result[1247:1235]);
small_alu1 sa96(clk, acc[1260:1248], secret[1260:1248], a_coeff, result[1260:1248]);
small_alu1 sa97(clk, acc[1273:1261], secret[1273:1261], a_coeff, result[1273:1261]);
small_alu1 sa98(clk, acc[1286:1274], secret[1286:1274], a_coeff, result[1286:1274]);
small_alu1 sa99(clk, acc[1299:1287], secret[1299:1287], a_coeff, result[1299:1287]);
small_alu1 sa100(clk, acc[1312:1300], secret[1312:1300], a_coeff, result[1312:1300]);
small_alu1 sa101(clk, acc[1325:1313], secret[1325:1313], a_coeff, result[1325:1313]);
small_alu1 sa102(clk, acc[1338:1326], secret[1338:1326], a_coeff, result[1338:1326]);
small_alu1 sa103(clk, acc[1351:1339], secret[1351:1339], a_coeff, result[1351:1339]);
small_alu1 sa104(clk, acc[1364:1352], secret[1364:1352], a_coeff, result[1364:1352]);
small_alu1 sa105(clk, acc[1377:1365], secret[1377:1365], a_coeff, result[1377:1365]);
small_alu1 sa106(clk, acc[1390:1378], secret[1390:1378], a_coeff, result[1390:1378]);
small_alu1 sa107(clk, acc[1403:1391], secret[1403:1391], a_coeff, result[1403:1391]);
small_alu1 sa108(clk, acc[1416:1404], secret[1416:1404], a_coeff, result[1416:1404]);
small_alu1 sa109(clk, acc[1429:1417], secret[1429:1417], a_coeff, result[1429:1417]);
small_alu1 sa110(clk, acc[1442:1430], secret[1442:1430], a_coeff, result[1442:1430]);
small_alu1 sa111(clk, acc[1455:1443], secret[1455:1443], a_coeff, result[1455:1443]);
small_alu1 sa112(clk, acc[1468:1456], secret[1468:1456], a_coeff, result[1468:1456]);
small_alu1 sa113(clk, acc[1481:1469], secret[1481:1469], a_coeff, result[1481:1469]);
small_alu1 sa114(clk, acc[1494:1482], secret[1494:1482], a_coeff, result[1494:1482]);
small_alu1 sa115(clk, acc[1507:1495], secret[1507:1495], a_coeff, result[1507:1495]);
small_alu1 sa116(clk, acc[1520:1508], secret[1520:1508], a_coeff, result[1520:1508]);
small_alu1 sa117(clk, acc[1533:1521], secret[1533:1521], a_coeff, result[1533:1521]);
small_alu1 sa118(clk, acc[1546:1534], secret[1546:1534], a_coeff, result[1546:1534]);
small_alu1 sa119(clk, acc[1559:1547], secret[1559:1547], a_coeff, result[1559:1547]);
small_alu1 sa120(clk, acc[1572:1560], secret[1572:1560], a_coeff, result[1572:1560]);
small_alu1 sa121(clk, acc[1585:1573], secret[1585:1573], a_coeff, result[1585:1573]);
small_alu1 sa122(clk, acc[1598:1586], secret[1598:1586], a_coeff, result[1598:1586]);
small_alu1 sa123(clk, acc[1611:1599], secret[1611:1599], a_coeff, result[1611:1599]);
small_alu1 sa124(clk, acc[1624:1612], secret[1624:1612], a_coeff, result[1624:1612]);
small_alu1 sa125(clk, acc[1637:1625], secret[1637:1625], a_coeff, result[1637:1625]);
small_alu1 sa126(clk, acc[1650:1638], secret[1650:1638], a_coeff, result[1650:1638]);
small_alu1 sa127(clk, acc[1663:1651], secret[1663:1651], a_coeff, result[1663:1651]);
small_alu1 sa128(clk, acc[1676:1664], secret[1676:1664], a_coeff, result[1676:1664]);
small_alu1 sa129(clk, acc[1689:1677], secret[1689:1677], a_coeff, result[1689:1677]);
small_alu1 sa130(clk, acc[1702:1690], secret[1702:1690], a_coeff, result[1702:1690]);
small_alu1 sa131(clk, acc[1715:1703], secret[1715:1703], a_coeff, result[1715:1703]);
small_alu1 sa132(clk, acc[1728:1716], secret[1728:1716], a_coeff, result[1728:1716]);
small_alu1 sa133(clk, acc[1741:1729], secret[1741:1729], a_coeff, result[1741:1729]);
small_alu1 sa134(clk, acc[1754:1742], secret[1754:1742], a_coeff, result[1754:1742]);
small_alu1 sa135(clk, acc[1767:1755], secret[1767:1755], a_coeff, result[1767:1755]);
small_alu1 sa136(clk, acc[1780:1768], secret[1780:1768], a_coeff, result[1780:1768]);
small_alu1 sa137(clk, acc[1793:1781], secret[1793:1781], a_coeff, result[1793:1781]);
small_alu1 sa138(clk, acc[1806:1794], secret[1806:1794], a_coeff, result[1806:1794]);
small_alu1 sa139(clk, acc[1819:1807], secret[1819:1807], a_coeff, result[1819:1807]);
small_alu1 sa140(clk, acc[1832:1820], secret[1832:1820], a_coeff, result[1832:1820]);
small_alu1 sa141(clk, acc[1845:1833], secret[1845:1833], a_coeff, result[1845:1833]);
small_alu1 sa142(clk, acc[1858:1846], secret[1858:1846], a_coeff, result[1858:1846]);
small_alu1 sa143(clk, acc[1871:1859], secret[1871:1859], a_coeff, result[1871:1859]);
small_alu1 sa144(clk, acc[1884:1872], secret[1884:1872], a_coeff, result[1884:1872]);
small_alu1 sa145(clk, acc[1897:1885], secret[1897:1885], a_coeff, result[1897:1885]);
small_alu1 sa146(clk, acc[1910:1898], secret[1910:1898], a_coeff, result[1910:1898]);
small_alu1 sa147(clk, acc[1923:1911], secret[1923:1911], a_coeff, result[1923:1911]);
small_alu1 sa148(clk, acc[1936:1924], secret[1936:1924], a_coeff, result[1936:1924]);
small_alu1 sa149(clk, acc[1949:1937], secret[1949:1937], a_coeff, result[1949:1937]);
small_alu1 sa150(clk, acc[1962:1950], secret[1962:1950], a_coeff, result[1962:1950]);
small_alu1 sa151(clk, acc[1975:1963], secret[1975:1963], a_coeff, result[1975:1963]);
small_alu1 sa152(clk, acc[1988:1976], secret[1988:1976], a_coeff, result[1988:1976]);
small_alu1 sa153(clk, acc[2001:1989], secret[2001:1989], a_coeff, result[2001:1989]);
small_alu1 sa154(clk, acc[2014:2002], secret[2014:2002], a_coeff, result[2014:2002]);
small_alu1 sa155(clk, acc[2027:2015], secret[2027:2015], a_coeff, result[2027:2015]);
small_alu1 sa156(clk, acc[2040:2028], secret[2040:2028], a_coeff, result[2040:2028]);
small_alu1 sa157(clk, acc[2053:2041], secret[2053:2041], a_coeff, result[2053:2041]);
small_alu1 sa158(clk, acc[2066:2054], secret[2066:2054], a_coeff, result[2066:2054]);
small_alu1 sa159(clk, acc[2079:2067], secret[2079:2067], a_coeff, result[2079:2067]);
small_alu1 sa160(clk, acc[2092:2080], secret[2092:2080], a_coeff, result[2092:2080]);
small_alu1 sa161(clk, acc[2105:2093], secret[2105:2093], a_coeff, result[2105:2093]);
small_alu1 sa162(clk, acc[2118:2106], secret[2118:2106], a_coeff, result[2118:2106]);
small_alu1 sa163(clk, acc[2131:2119], secret[2131:2119], a_coeff, result[2131:2119]);
small_alu1 sa164(clk, acc[2144:2132], secret[2144:2132], a_coeff, result[2144:2132]);
small_alu1 sa165(clk, acc[2157:2145], secret[2157:2145], a_coeff, result[2157:2145]);
small_alu1 sa166(clk, acc[2170:2158], secret[2170:2158], a_coeff, result[2170:2158]);
small_alu1 sa167(clk, acc[2183:2171], secret[2183:2171], a_coeff, result[2183:2171]);
small_alu1 sa168(clk, acc[2196:2184], secret[2196:2184], a_coeff, result[2196:2184]);
small_alu1 sa169(clk, acc[2209:2197], secret[2209:2197], a_coeff, result[2209:2197]);
small_alu1 sa170(clk, acc[2222:2210], secret[2222:2210], a_coeff, result[2222:2210]);
small_alu1 sa171(clk, acc[2235:2223], secret[2235:2223], a_coeff, result[2235:2223]);
small_alu1 sa172(clk, acc[2248:2236], secret[2248:2236], a_coeff, result[2248:2236]);
small_alu1 sa173(clk, acc[2261:2249], secret[2261:2249], a_coeff, result[2261:2249]);
small_alu1 sa174(clk, acc[2274:2262], secret[2274:2262], a_coeff, result[2274:2262]);
small_alu1 sa175(clk, acc[2287:2275], secret[2287:2275], a_coeff, result[2287:2275]);
small_alu1 sa176(clk, acc[2300:2288], secret[2300:2288], a_coeff, result[2300:2288]);
small_alu1 sa177(clk, acc[2313:2301], secret[2313:2301], a_coeff, result[2313:2301]);
small_alu1 sa178(clk, acc[2326:2314], secret[2326:2314], a_coeff, result[2326:2314]);
small_alu1 sa179(clk, acc[2339:2327], secret[2339:2327], a_coeff, result[2339:2327]);
small_alu1 sa180(clk, acc[2352:2340], secret[2352:2340], a_coeff, result[2352:2340]);
small_alu1 sa181(clk, acc[2365:2353], secret[2365:2353], a_coeff, result[2365:2353]);
small_alu1 sa182(clk, acc[2378:2366], secret[2378:2366], a_coeff, result[2378:2366]);
small_alu1 sa183(clk, acc[2391:2379], secret[2391:2379], a_coeff, result[2391:2379]);
small_alu1 sa184(clk, acc[2404:2392], secret[2404:2392], a_coeff, result[2404:2392]);
small_alu1 sa185(clk, acc[2417:2405], secret[2417:2405], a_coeff, result[2417:2405]);
small_alu1 sa186(clk, acc[2430:2418], secret[2430:2418], a_coeff, result[2430:2418]);
small_alu1 sa187(clk, acc[2443:2431], secret[2443:2431], a_coeff, result[2443:2431]);
small_alu1 sa188(clk, acc[2456:2444], secret[2456:2444], a_coeff, result[2456:2444]);
small_alu1 sa189(clk, acc[2469:2457], secret[2469:2457], a_coeff, result[2469:2457]);
small_alu1 sa190(clk, acc[2482:2470], secret[2482:2470], a_coeff, result[2482:2470]);
small_alu1 sa191(clk, acc[2495:2483], secret[2495:2483], a_coeff, result[2495:2483]);
small_alu1 sa192(clk, acc[2508:2496], secret[2508:2496], a_coeff, result[2508:2496]);
small_alu1 sa193(clk, acc[2521:2509], secret[2521:2509], a_coeff, result[2521:2509]);
small_alu1 sa194(clk, acc[2534:2522], secret[2534:2522], a_coeff, result[2534:2522]);
small_alu1 sa195(clk, acc[2547:2535], secret[2547:2535], a_coeff, result[2547:2535]);
small_alu1 sa196(clk, acc[2560:2548], secret[2560:2548], a_coeff, result[2560:2548]);
small_alu1 sa197(clk, acc[2573:2561], secret[2573:2561], a_coeff, result[2573:2561]);
small_alu1 sa198(clk, acc[2586:2574], secret[2586:2574], a_coeff, result[2586:2574]);
small_alu1 sa199(clk, acc[2599:2587], secret[2599:2587], a_coeff, result[2599:2587]);
small_alu1 sa200(clk, acc[2612:2600], secret[2612:2600], a_coeff, result[2612:2600]);
small_alu1 sa201(clk, acc[2625:2613], secret[2625:2613], a_coeff, result[2625:2613]);
small_alu1 sa202(clk, acc[2638:2626], secret[2638:2626], a_coeff, result[2638:2626]);
small_alu1 sa203(clk, acc[2651:2639], secret[2651:2639], a_coeff, result[2651:2639]);
small_alu1 sa204(clk, acc[2664:2652], secret[2664:2652], a_coeff, result[2664:2652]);
small_alu1 sa205(clk, acc[2677:2665], secret[2677:2665], a_coeff, result[2677:2665]);
small_alu1 sa206(clk, acc[2690:2678], secret[2690:2678], a_coeff, result[2690:2678]);
small_alu1 sa207(clk, acc[2703:2691], secret[2703:2691], a_coeff, result[2703:2691]);
small_alu1 sa208(clk, acc[2716:2704], secret[2716:2704], a_coeff, result[2716:2704]);
small_alu1 sa209(clk, acc[2729:2717], secret[2729:2717], a_coeff, result[2729:2717]);
small_alu1 sa210(clk, acc[2742:2730], secret[2742:2730], a_coeff, result[2742:2730]);
small_alu1 sa211(clk, acc[2755:2743], secret[2755:2743], a_coeff, result[2755:2743]);
small_alu1 sa212(clk, acc[2768:2756], secret[2768:2756], a_coeff, result[2768:2756]);
small_alu1 sa213(clk, acc[2781:2769], secret[2781:2769], a_coeff, result[2781:2769]);
small_alu1 sa214(clk, acc[2794:2782], secret[2794:2782], a_coeff, result[2794:2782]);
small_alu1 sa215(clk, acc[2807:2795], secret[2807:2795], a_coeff, result[2807:2795]);
small_alu1 sa216(clk, acc[2820:2808], secret[2820:2808], a_coeff, result[2820:2808]);
small_alu1 sa217(clk, acc[2833:2821], secret[2833:2821], a_coeff, result[2833:2821]);
small_alu1 sa218(clk, acc[2846:2834], secret[2846:2834], a_coeff, result[2846:2834]);
small_alu1 sa219(clk, acc[2859:2847], secret[2859:2847], a_coeff, result[2859:2847]);
small_alu1 sa220(clk, acc[2872:2860], secret[2872:2860], a_coeff, result[2872:2860]);
small_alu1 sa221(clk, acc[2885:2873], secret[2885:2873], a_coeff, result[2885:2873]);
small_alu1 sa222(clk, acc[2898:2886], secret[2898:2886], a_coeff, result[2898:2886]);
small_alu1 sa223(clk, acc[2911:2899], secret[2911:2899], a_coeff, result[2911:2899]);
small_alu1 sa224(clk, acc[2924:2912], secret[2924:2912], a_coeff, result[2924:2912]);
small_alu1 sa225(clk, acc[2937:2925], secret[2937:2925], a_coeff, result[2937:2925]);
small_alu1 sa226(clk, acc[2950:2938], secret[2950:2938], a_coeff, result[2950:2938]);
small_alu1 sa227(clk, acc[2963:2951], secret[2963:2951], a_coeff, result[2963:2951]);
small_alu1 sa228(clk, acc[2976:2964], secret[2976:2964], a_coeff, result[2976:2964]);
small_alu1 sa229(clk, acc[2989:2977], secret[2989:2977], a_coeff, result[2989:2977]);
small_alu1 sa230(clk, acc[3002:2990], secret[3002:2990], a_coeff, result[3002:2990]);
small_alu1 sa231(clk, acc[3015:3003], secret[3015:3003], a_coeff, result[3015:3003]);
small_alu1 sa232(clk, acc[3028:3016], secret[3028:3016], a_coeff, result[3028:3016]);
small_alu1 sa233(clk, acc[3041:3029], secret[3041:3029], a_coeff, result[3041:3029]);
small_alu1 sa234(clk, acc[3054:3042], secret[3054:3042], a_coeff, result[3054:3042]);
small_alu1 sa235(clk, acc[3067:3055], secret[3067:3055], a_coeff, result[3067:3055]);
small_alu1 sa236(clk, acc[3080:3068], secret[3080:3068], a_coeff, result[3080:3068]);
small_alu1 sa237(clk, acc[3093:3081], secret[3093:3081], a_coeff, result[3093:3081]);
small_alu1 sa238(clk, acc[3106:3094], secret[3106:3094], a_coeff, result[3106:3094]);
small_alu1 sa239(clk, acc[3119:3107], secret[3119:3107], a_coeff, result[3119:3107]);
small_alu1 sa240(clk, acc[3132:3120], secret[3132:3120], a_coeff, result[3132:3120]);
small_alu1 sa241(clk, acc[3145:3133], secret[3145:3133], a_coeff, result[3145:3133]);
small_alu1 sa242(clk, acc[3158:3146], secret[3158:3146], a_coeff, result[3158:3146]);
small_alu1 sa243(clk, acc[3171:3159], secret[3171:3159], a_coeff, result[3171:3159]);
small_alu1 sa244(clk, acc[3184:3172], secret[3184:3172], a_coeff, result[3184:3172]);
small_alu1 sa245(clk, acc[3197:3185], secret[3197:3185], a_coeff, result[3197:3185]);
small_alu1 sa246(clk, acc[3210:3198], secret[3210:3198], a_coeff, result[3210:3198]);
small_alu1 sa247(clk, acc[3223:3211], secret[3223:3211], a_coeff, result[3223:3211]);
small_alu1 sa248(clk, acc[3236:3224], secret[3236:3224], a_coeff, result[3236:3224]);
small_alu1 sa249(clk, acc[3249:3237], secret[3249:3237], a_coeff, result[3249:3237]);
small_alu1 sa250(clk, acc[3262:3250], secret[3262:3250], a_coeff, result[3262:3250]);
small_alu1 sa251(clk, acc[3275:3263], secret[3275:3263], a_coeff, result[3275:3263]);
small_alu1 sa252(clk, acc[3288:3276], secret[3288:3276], a_coeff, result[3288:3276]);
small_alu1 sa253(clk, acc[3301:3289], secret[3301:3289], a_coeff, result[3301:3289]);
small_alu1 sa254(clk, acc[3314:3302], secret[3314:3302], a_coeff, result[3314:3302]);
small_alu1 sa255(clk, acc[3327:3315], secret[3327:3315], a_coeff, result[3327:3315]);

endmodule
