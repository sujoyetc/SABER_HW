module s_rom(clk, s_address, s_vec_64);
input clk;
input [6:0] s_address;
output reg [63:0] s_vec_64;

wire [63:0] s_vec_64_wire;

/*
assign s_vec_64_wire =	
						(s_address==7'd0) ? 64'b1010000110011001001100100011001010100011100110111011101100110011:
            (s_address==7'd1) ? 64'b0001000000011001000100110010001100000010000010100010000110110001:
            (s_address==7'd2) ? 64'b1011101010101010000110100001000000001001000010011011001110111001:
            (s_address==7'd3) ? 64'b0001001000000011000010100001001000011001000100011010101010011010:
            (s_address==7'd4) ? 64'b0001001000000010001000000011101000000011100110010001001110010011:
            (s_address==7'd5) ? 64'b0001001000011001000000000010100100110011000100010000100100001010:
            (s_address==7'd6) ? 64'b1001100100000011100100011010001100100011100110100010000000000010:
            (s_address==7'd7) ? 64'b0001000010100010100100000001000100100001000100010001001100100011:
            (s_address==7'd8) ? 64'b0010000110111011001010100011101100101001001100111011000100101001:
            (s_address==7'd9) ? 64'b0000101110100011101010010011101000010011101100101010000110011011:
            (s_address==7'd10) ? 64'b0010101110111011101110111011001010101010100110011011101100110010:
            (s_address==7'd11) ? 64'b1010001110110001000010110010000110100010101000111010100110011011:
            (s_address==7'd12) ? 64'b0001000010011011000010011001101100100010001000011001101110111010:
            (s_address==7'd13) ? 64'b0010001010111010000010100010000100110000001110011011001000010011:
            (s_address==7'd14) ? 64'b1010100100010000000000110001000110100011001100001011101100111001:
            (s_address==7'd15) ? 64'b1010101110011011001010100001001010110010000000011001100110010011: 64'd0;
*/

assign s_vec_64_wire =	
						(s_address==7'd0) ? 64'b10001010110001101010010001000110011001000110001000100010000001:
						(s_address==7'd1) ? 64'b1010101110000010100100001001001010110011000100000010101000001011:
						(s_address==7'd2) ? 64'b1011001110001011001000100010000010110000100100101011001000101011:
						(s_address==7'd3) ? 64'b100000111010001110001000001110001010001000010000000110111000:
						(s_address==7'd4) ? 64'b1101000001000000010110001000000010000001100110001000110110000:
						(s_address==7'd5) ? 64'b1001110001000101010001010000100010000100110001000101000011010:
						(s_address==7'd6) ? 64'b1011001000000011100100110011001110011000100000011001100000110001:
						(s_address==7'd7) ? 64'b1001001000010011000110001010100110110010000010010001101000100000:
						(s_address==7'd8) ? 64'b11101100001010000100111000001010000000000100000000100010100010:
						(s_address==7'd9) ? 64'b10100110111010101000100000101100001010101100101000101100010000:
						(s_address==7'd10) ? 64'b1011001110001000000000011011001100011001101100011001000000111011:
						(s_address==7'd11) ? 64'b1011000110101000101000010010000100010011100110001011101110110001:
						(s_address==7'd12) ? 64'b1010001010100010100010110000001100011010001110010001100100111001:
						(s_address==7'd13) ? 64'b1000100001001001100100000001010000000101010000010101110111011:
						(s_address==7'd14) ? 64'b11000110100000100100010000000110110010100010101011101000000001:
						(s_address==7'd15) ? 64'b11000110110011000000111000101100111011101010001001000010000001:64'b0;

always @(posedge clk)
	s_vec_64 <= s_vec_64_wire;
	
endmodule
