module s_rom(clk, s_address, s_vec_64);
input clk;
input [6:0] s_address;
output reg [63:0] s_vec_64;

wire [63:0] s_vec_64_wire;

assign s_vec_64_wire =	
						(s_address==7'd0) ? 64'b1010000110011001001100100011001010100011100110111011101100110011:
            (s_address==7'd1) ? 64'b0001000000011001000100110010001100000010000010100010000110110001:
            (s_address==7'd2) ? 64'b1011101010101010000110100001000000001001000010011011001110111001:
            (s_address==7'd3) ? 64'b0001001000000011000010100001001000011001000100011010101010011010:
            (s_address==7'd4) ? 64'b0001001000000010001000000011101000000011100110010001001110010011:
            (s_address==7'd5) ? 64'b0001001000011001000000000010100100110011000100010000100100001010:
            (s_address==7'd6) ? 64'b1001100100000011100100011010001100100011100110100010000000000010:
            (s_address==7'd7) ? 64'b0001000010100010100100000001000100100001000100010001001100100011:
            (s_address==7'd8) ? 64'b0010000110111011001010100011101100101001001100111011000100101001:
            (s_address==7'd9) ? 64'b0000101110100011101010010011101000010011101100101010000110011011:
            (s_address==7'd10) ? 64'b0010101110111011101110111011001010101010100110011011101100110010:
            (s_address==7'd11) ? 64'b1010001110110001000010110010000110100010101000111010100110011011:
            (s_address==7'd12) ? 64'b0001000010011011000010011001101100100010001000011001101110111010:
            (s_address==7'd13) ? 64'b0010001010111010000010100010000100110000001110011011001000010011:
            (s_address==7'd14) ? 64'b1010100100010000000000110001000110100011001100001011101100111001:
            (s_address==7'd15) ? 64'b1010101110011011001010100001001010110010000000011001100110010011: 64'd0;

always @(posedge clk)
	s_vec_64 <= s_vec_64_wire;
	
endmodule
