module pol_rom(clk, bram_address_relative, pol_64bit_in);
input clk;
input [6:0] bram_address_relative;
output reg [63:0] pol_64bit_in;

wire [63:0] pol_64bit_in_wire;
assign pol_64bit_in_wire = 	
						(bram_address_relative==7'd0) ?  64'b1110110100111110100000100001100010001001010111011000101001010000:
            (bram_address_relative==7'd1) ?  64'b1001011010111100011101010111011100000011111100101000010000000100:
            (bram_address_relative==7'd2) ?  64'b0001101100101110000011101110100110100010100100101100000000110000:
            (bram_address_relative==7'd3) ?  64'b0010001010100110101011000000100111110001110101101101100010010100:
            (bram_address_relative==7'd4) ?  64'b1001111000111000111010101001000001110100010100011000100111110001:
            (bram_address_relative==7'd5) ?  64'b0100001000010100010000110011000100011010000101011110110101000101:
            (bram_address_relative==7'd6) ?  64'b1110000000110010000011011110100100110101110110111011010001010111:
            (bram_address_relative==7'd7) ?  64'b1001001101100110001100001010001100111101001011101000011001110110:
            (bram_address_relative==7'd8) ?  64'b0000000110100011100001010111011101100111101110111100001001101011:
            (bram_address_relative==7'd9) ?  64'b1111011101101111111101011010100110000000000101110011001110101100:
            (bram_address_relative==7'd10) ?  64'b1010111110100101001010001000101110111010000111100101100000100111:
            (bram_address_relative==7'd11) ?  64'b0001101011100000110011110011101001100010000010011100010011101110:
            (bram_address_relative==7'd12) ?  64'b0001111010110111001110010000001000000010110010110010100111001010:
            (bram_address_relative==7'd13) ?  64'b0100101110000110101010011111011010011111111000110001101001001000:
            (bram_address_relative==7'd14) ?  64'b0111001001010111110111010000110001011100100011001000000010101110:
            (bram_address_relative==7'd15) ?  64'b1101101000011000100111111111011000110111000000110001001110011010:
            (bram_address_relative==7'd16) ?  64'b0000100110100011110000111011010010111001000100101011111100101001:
            (bram_address_relative==7'd17) ?  64'b1101111000111110010111000001000100001111100101011001010010001011:
            (bram_address_relative==7'd18) ?  64'b0111110011011001000111001000001111010101101000001010010011100111:
            (bram_address_relative==7'd19) ?  64'b0110111111111011110000101100001111110000110100000110010100001101:
            (bram_address_relative==7'd20) ?  64'b1011010111111111100100100001101111010100000010110111000101001010:
            (bram_address_relative==7'd21) ?  64'b1110111110111111011010110100001111010010000111101111110110001001:
            (bram_address_relative==7'd22) ?  64'b0101111101001000010100000001001110110100101100101000010100101111:
            (bram_address_relative==7'd23) ?  64'b0100100100011010011000100100001010110010111011010111101000010011:
            (bram_address_relative==7'd24) ?  64'b1001000100011111010101011000100101100000010110100010110110110010:
            (bram_address_relative==7'd25) ?  64'b1100011111111100101111011101000001110010001001100111001011000001:
            (bram_address_relative==7'd26) ?  64'b0010010111100101100001010111000001011010101000101010111011010100:
            (bram_address_relative==7'd27) ?  64'b1010000101100110001001111101100011110010011111110000111001011001:
            (bram_address_relative==7'd28) ?  64'b0110000000010100001010001010110110101000001110110011111110100110:
            (bram_address_relative==7'd29) ?  64'b1110111010100101000011101101111001011001110111010111100000001111:
            (bram_address_relative==7'd30) ?  64'b0010010001011100011001100010000111000011110000111100001111001110:
            (bram_address_relative==7'd31) ?  64'b0111100110011110101010001100010001111011100000000110110110111001:
            (bram_address_relative==7'd32) ?  64'b1101011010100101010101110000101111110001111011101001100000100000:
            (bram_address_relative==7'd33) ?  64'b1111011000011110111100111000110011000000011001110011001100010100:
            (bram_address_relative==7'd34) ?  64'b1011010110101101011101110101111110110111011101000000011100000101:
            (bram_address_relative==7'd35) ?  64'b0101100010110000011011101101111001110010010000100011000001100000:
            (bram_address_relative==7'd36) ?  64'b0110001100011110110011000101110001111010100110011011010110111001:
            (bram_address_relative==7'd37) ?  64'b0110111100110100000100010110100011010010111110101100001100010000:
            (bram_address_relative==7'd38) ?  64'b0110100011110111011110010001011000110111000000111100111101101101:
            (bram_address_relative==7'd39) ?  64'b0100001100001111100010001000000011000110110011010100010010101001:
            (bram_address_relative==7'd40) ?  64'b1010111010110001000101011110101100101101010110111011111000010100:
            (bram_address_relative==7'd41) ?  64'b0111100011010110001110110110001111110010100011011000011100001111:
            (bram_address_relative==7'd42) ?  64'b1111101110101001100111000110111011001000101000011000001010110110:
            (bram_address_relative==7'd43) ?  64'b1010101001001111110011001011011110111011011110011000011011011111:
            (bram_address_relative==7'd44) ?  64'b0101101101110111010000000000111011110111101001100100001011100000:
            (bram_address_relative==7'd45) ?  64'b1000111001110111101011010001010111100010101101100001111000000100:
            (bram_address_relative==7'd46) ?  64'b0001000100111010001001101011111111101111011001000100010011111111:
            (bram_address_relative==7'd47) ?  64'b0110100111111101010101010110111001101110111101000000100110000100:
            (bram_address_relative==7'd48) ?  64'b1000100110010010110010000100001101011110100010111110010110010010:
            (bram_address_relative==7'd49) ?  64'b1011101010010000111011101000000101001111110011101101110010110110:
            (bram_address_relative==7'd50) ?  64'b1001110010101000111001010010001111101011100011100001001110110110:
            (bram_address_relative==7'd51) ?  64'b1011011001010101000110000001101101011011011101010101110000100010: 
						64'd0;
						
		always @(posedge clk)
			pol_64bit_in <= pol_64bit_in_wire;
			
endmodule
			
		